magic
tech sky130A
magscale 1 2
timestamp 1769042447
<< locali >>
rect 192 1960 425 2040
rect -96 -200 96 200
rect 1056 -200 1248 152
rect -400 -208 1600 -200
rect -400 -388 294 -208
rect 474 -388 1600 -208
rect -400 -400 1600 -388
<< viali >>
rect 294 -388 474 -208
<< metal1 >>
rect 160 544 224 3907
rect 160 360 224 440
rect 288 -208 480 3806
rect 673 3240 1200 3430
rect 1000 2632 1200 3240
rect 672 2440 1200 2632
rect 1000 1560 1200 2440
rect 672 1368 1200 1560
rect 1000 760 1200 1368
rect 672 568 1200 760
rect 1000 400 1200 568
rect 672 40 864 120
rect 288 -388 294 -208
rect 474 -388 480 -208
rect 288 -400 480 -388
use JNWATR_NCH_4C5F0  xo0<0> ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 0
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo0<1>
timestamp 1740610800
transform 1 0 0 0 1 800
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1
timestamp 1740610800
transform 1 0 0 0 1 1600
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo2<0>
timestamp 1740610800
transform 1 0 0 0 1 2400
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo2<1>
timestamp 1740610800
transform 1 0 0 0 1 3200
box -184 -128 1336 928
<< labels >>
flabel metal1 s 672 40 864 120 0 FreeSans 400 0 0 0 IBNS_20U
port 1 nsew signal bidirectional
flabel metal1 s 288 600 480 680 0 FreeSans 400 0 0 0 VSS
port 2 nsew ground bidirectional
flabel metal1 s 160 360 224 440 0 FreeSans 400 0 0 0 IBPS_5U
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 4000
<< end >>
